`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:31:21 01/05/2019 
// Design Name: 
// Module Name:    IsHit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module IsHit(
input wire clk,
	input wire  [9:0] ebi_x,
	input wire  [8:0] ebi_y,
	input wire  [9:0] mi_x,
	input wire  [8:0] mi_y,
	output wire check
    );
	 reg [9:0] e_xm;
	 reg [8:0] e_ym;
	  
	 reg [9:0] m_x;
	 reg [8:0] m_y;
	 
	 reg in;
	 
	 integer k;
	 
	 always @(posedge clk) begin
		 e_xm<=ebi_x;
		 e_ym<=ebi_y;
		 	 
		 m_x<=mi_x+40;
		 m_y<=mi_y+41;
		 in = 0;
		 k = 30;
		 if(e_xm< m_x+38 && e_xm>m_x-38 && e_ym <m_y+38 && e_ym >m_y-38) begin//in the square
				if(e_ym<m_y) begin
					if(e_xm<m_x)begin
						k= m_x- e_xm + m_y- e_ym;
					end
					else begin
						k= e_xm-m_x + m_y- e_ym;
					end			
				end
				if(k<38) begin
					in = 1;
				end
		 end
	end
	
	assign check = in;
	 




endmodule
